Entity Laboratory1A is
end entity;

architecture sim of Laboratory1A is
begin

process is
begin
		
	report "Marco, Roldan L.";
	report "20101140787";
	report "BSCpE";
	wait;

end process;

end architecture;