Entity Laboratory1A is
end entity;

architecture sim of Laboratory1A is
begin

process is
begin
		
	report "Marco, Roldan L.";
	wait for 1000 ms;
	report "20101140787";
	wait for 1000 ms;
	report "BSCpE";
	wait;

end process;

end architecture;
